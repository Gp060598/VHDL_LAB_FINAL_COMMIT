// The mem_type should be converted into a class so that you can collect statistics of the instructions

typedef bit [15:0] uint16;
typedef uint16 mem_type;

class mem_class;
endclass
